module enums

pub enum Align {
	left
	center
	right
	justify
}
