module enums

pub enum Dock {
	top
	bottom
	left
	right
}
