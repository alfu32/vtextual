module geometry

import geometry { Point, Size }

pub struct Region {
pub:
	origin Point
	size   Size
}
