module main

fn main() {
	dump('Hello World!')
}
