module geometry

pub struct Spacing {
pub:
	horizontal int
	vertical   int
}
